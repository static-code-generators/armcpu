`define S_BIT 20

`define L_BIT 20
`define W_BIT 21
`define B_BIT 22
`define U_BIT 23
`define P_BIT 24
`define I_BIT 25

`define EQ 0000
`define NE 0001
`define CS 0010
`define CC 0011
`define MI 0100
`define PL 0101
`define VS 0110
`define VC 0111
`define HI 1000
`define LS 1001
`define GE 1010
`define LT 1011
`define GT 1100
`define LE 1101
`define AL 1110
