`define NULL 0
`define TEST_FILE_NAME "test/additest.x"

module tb_final;

    reg        clk;
    wire [1:0] we;
    wire [1:0] excpt;

    assign we[0] = 1'b0;
    assign we[1] = mem_write_en;

    arm_memory memauri
    (
        // Inputs
        .clk(clk),
        .addr1(inst_addr),
        .addr2(mem_addr),
        .data_in1(),
        .data_in2(mem_data_in),
        .we(we),
        .excpt(excpt),
        // Outputs
        .data_out1(inst),
        .data_out2(mem_data_out)
    );

    arm_core core
    (
        // Inputs
        .clk(clk),
        .rst(rst),
        .inst(inst),
        .mem_data_out(mem_data_out),
        // Outputs
        .halted(halted),
        .mem_addr(mem_addr),
        .inst_addr(inst_addr),
        .mem_data_in(mem_data_in)
        .mem_write_en(mem_write_en)
    );

    always #10 clk = ~clk;

    integer index;

    initial begin
        index = 0;
        clk = 0;
        rst = 1;
        text_file = $fopen(`TEST_FILE_NAME, "r");

        if (data_file == `NULL) begin
            $display("bad bad | text file handle was NULL");
            $finish;
        end
    end

    always @(negedge clk) begin
        scan_file = $fscanf(text_file, "%x\n", captured_data);
        if (!$feof(text_file)) begin
            $display("read from file: %x, trying to write to: %d",
            mem_data_in, index);
            //mem_write_en = 0; //not ready to write yet.
            mem_addr = index;
            mem_write_en = 1;
            index = index + 4;
        end
        else begin
            rst = 0;
            if (halted)
                #10 $finish;
        end
    end

endmodule
