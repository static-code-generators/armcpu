module barrel_shifter
(
    input      [31:0] inst;
    output reg [31:0] shifter_operand;
    output reg [31:0] shifter_carry;
);

// fill me up bby

endmodule
