`include "arm_defines.vh"

/*
 * Outputs valid signal depending on current status of CPSR
 */
module cond_decode
(
    // inputs
    input [31:0] inst, cpsr,
    // outputs
    output valid
);

    // Stuff in the cases here

endmodule
